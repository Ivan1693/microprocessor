library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom3216 is
    Port ( address : in std_logic_vector (4 downto 0);
           data : out  std_logic_vector (15 downto 0));
end rom3216;

architecture behavioral of rom3216 is
	type reg_grid is array (31 downto 0) of std_logic_vector(15 downto 0);
constant rom: reg_grid := (
"1000000000010010",
"0111000010101111",
"1000000000011000",
"1000000000010111",
"1000000000010110",
"1000000000010101",
"1000000000010100",
"1000000000011110",
"1000000000011101",
"1000000000011100",
"1000000000011011",
"1000000000011010",
"1000000000011001",
"0111000010101111",
"0111110110001111",
"0011100110001111",
"0011010010001101",
"0011000110100100",
"0110110000000101",
"0110100101000110",
"0010010011101111",
"0010000011001010",
"0100010000010101",
"0001111111000101",
"0001101111000101",
"0101010011000001",
"0000110011000001",
"0001000011101101",
"0000100011101101",
"0100000000011011",
"0000010110000100",
"0000000100000011"
);
begin
	data <= rom(to_integer(unsigned(address)));
end architecture;