library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom3216 is
    Port ( address : in std_logic_vector (4 downto 0);
           data : out  std_logic_vector (15 downto 0));
end rom3216;

architecture behavioral of rom3216 is
	type reg_grid is array (31 downto 0) of std_logic_vector(15 downto 0);
constant rom: reg_grid := (
"1100000001000001",--Guarda 00001 en 00001
"0000000000100000",--Suma los valores en las direcciones 00001 y 00000
"1110000000111111",--Transfiere el valor en el acumulador a la direccion 00001
"1000000000010110",
"1000000000010101",
"1000000000010100",
"1000000000011110",
"1000000000011101",
"1000000000011100",
"1000000000011011",
"1000000000011010",
"1000000000011001",
"0111000010101111",
"0111110111101100",
"0011100110001111",
"0011010010001101",
"0011000110100100",
"0110110000000101",
"0110100101000110",
"0010010011101111",
"0010000011001010",
"1000000000000011",--0x0A salto 0x03
"1110000000111111",--0x09 mov(ACM,00001)
"0000110000000001",--0x08 00001++
"1110000001011111",--0x07 mov(ACM,00010)
"0000000001000001",--0x06 sum(00010,00001)
"1000000000000101",--0x05 kill
"1000000000000110",--0x04 Salta a 0x06
"0011000000000001",--0x03 Si 00001 > 00000
"1100000000000010",--0x02 Guarda 00000 en 00010
"1100000000000001",--0x01 Guarda 00000 en 00001
"1100000011000000" --0x00 Guarda 00011 en 00000
);
begin
	data <= rom(to_integer(unsigned(address)));
end architecture;