library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity rom3216 is
    Port ( address : in std_logic_vector (4 downto 0);
           data : out  std_logic_vector (15 downto 0));
end rom3216;

architecture behavioral of rom3216 is
	type reg_grid is array (31 downto 0) of std_logic_vector(15 downto 0);
	constant rom: reg_grid := (
		--Zaid
		"0000000000000000",
		"1000000000000001",
		"0000000000000010",
		"0000000000000011",
		"0000000000000100",
		"0000000000000101",
		"0000000000000110",
		"0000000000000111",
		"0000000000001000",
		"0000000000001001",
		"1000000000011110",

		--Ramses
		"0011010001100110",
		"0011000101000101",
		"0001001010100000",
		"0001000010100000",
		"0001100000001110",
		"0001100000011110",
		"0000110000001111",
		"0000110000011110",
		"0000011101000010",
		"0000000101010010",

		--Ivan
		"0000000011101000",
		"0011110000000101",
		"0001110011100101",
		"0001100011100101",
		"0001010011000001",
		"0000110011000001",
		"0101000000001101",
		"0100100000001101",
		"0100000000011011",
		"0000010110000100",
		"0000000100000011");
begin
	data <= rom(to_integer(unsigned(address)));
end architecture;

