library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity rom3216 is
    Port ( address : in STD_LOGIC_VECTOR (4 downto 0);
           data : out  STD_LOGIC_VECTOR (15 downto 0));
end rom3216;

architecture Behavioral of rom3216 is
	type reg_grid is array (31 downto 0) of std_logic_vector(15 downto 0);
	constant rom: reg_grid := (
		"0000000000000000","0000000000000001","0000000000000010","0000000000000011",
		"0000000000000100","0000000000000101","0000000000000110","0000000000000111",
		"0000000000001000","0000000000001001","0000000000001010","0000000000001011",
		"0000000000001100","0000000000011101","0000000000001110","0000000000001111",
		"0000000000010000","0000000000010001","0000000000010010","0000000000010011",
		"0000000000010100","0000000000010101","0000000000010110","0000000000010111",
		"0000000000011000","0000000000011001","0000000000011010","0000000000011011",
		"0000000000011100","0000000000011101","0000000000011110","0000000000011111");
begin
	data <= rom(to_integer(unsigned(address)));
end Behavioral;

